`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:03:58 09/13/2020 
// Design Name: 
// Module Name:    eight_bit_cmparator 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module eight_bit_comparator(
    input [0:7] a,
    input [0:7] b,
    output G,
    output Eq,
    output L
    );
	
	one_bit_comparator c0();

endmodule
